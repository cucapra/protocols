module identity_d0 (
    input              clk,
    input       a,
    input       b,
    output      s1,
    output      s2
);
    assign s1 = a;
    assign s2 = b;
endmodule
